rustlightProbe_inst : rustlightProbe PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
