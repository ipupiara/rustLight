inputProbe_inst : inputProbe PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
