clkCtrlOut_inst : clkCtrlOut PORT MAP (
		inclk	 => inclk_sig,
		outclk	 => outclk_sig
	);
