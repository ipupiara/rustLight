triacDriverProbe_inst : triacDriverProbe PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
