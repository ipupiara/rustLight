demuxInputChecker_inst : demuxInputChecker PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
