controllerInputChecker_inst : controllerInputChecker PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
