rustLightCompare_1_inst : rustLightCompare_1 PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
